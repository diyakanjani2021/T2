<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>37.7991,72.5626,553.592,-182.384</PageViewport>
<gate>
<ID>390</ID>
<type>GA_LED</type>
<position>530.5,-83.5</position>
<input>
<ID>N_in0</ID>203 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>391</ID>
<type>AA_LABEL</type>
<position>522.5,-40</position>
<gparam>LABEL_TEXT FULL ADDER WITH NAND</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>32,-19</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>24,-18</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>24,-20</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>38,-19</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>31,-14.5</position>
<gparam>LABEL_TEXT AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>21,-17.5</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>21,-19.5</position>
<gparam>LABEL_TEXT i/p b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>42,-18.5</position>
<gparam>LABEL_TEXT y = ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>29,-22</position>
<gparam>LABEL_TEXT a b y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>29,-23.5</position>
<gparam>LABEL_TEXT 0 0 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>29.5,-26</position>
<gparam>LABEL_TEXT OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>32.5,-31</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>24,-30</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>24,-32</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>38.5,-31</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>20.5,-29.5</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>20.5,-31.5</position>
<gparam>LABEL_TEXT i/p b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>43,-30.5</position>
<gparam>LABEL_TEXT y = a+b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>30,-35.5</position>
<gparam>LABEL_TEXT NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>BE_NOR2</type>
<position>33,-40</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>24,-39</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>24,-41</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>39,-40</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>43.5,-39.5</position>
<gparam>LABEL_TEXT y = a+b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>20.5,-38.5</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>20.5,-40.5</position>
<gparam>LABEL_TEXT i/p b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>45,-37</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>30.5,-44.5</position>
<gparam>LABEL_TEXT NAND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>BA_NAND2</type>
<position>33.5,-49.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_TOGGLE</type>
<position>24.5,-48.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>24.5,-50.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>55,-18.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>39.5,-49.5</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>21,-48</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>21,-50</position>
<gparam>LABEL_TEXT i/p b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>43.5,-49</position>
<gparam>LABEL_TEXT y = ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>45,-46.5</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>62,-14.5</position>
<gparam>LABEL_TEXT NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_INVERTER</type>
<position>61.5,-18.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>67,-18.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>51.5,-18</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>71,-18</position>
<gparam>LABEL_TEXT y = a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>72.5,-15.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>62,-23</position>
<gparam>LABEL_TEXT XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AI_XOR2</type>
<position>65.5,-28.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>58,-27.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>58,-29.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>70.5,-28.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>54.5,-27.5</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>54.5,-29.5</position>
<gparam>LABEL_TEXT i/p b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>77,-28</position>
<gparam>LABEL_TEXT y = ab + ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>76,-25.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>81,-25.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>63,-33</position>
<gparam>LABEL_TEXT XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AO_XNOR2</type>
<position>66.5,-38</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>59,-37</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>59,-39</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>71.5,-38</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>56,-37</position>
<gparam>LABEL_TEXT i/p a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>56,-38.5</position>
<gparam>LABEL_TEXT i/p b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>77.5,-37.5</position>
<gparam>LABEL_TEXT y = ab + ab</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>81,-35</position>
<gparam>LABEL_TEXT __</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>121.5,-12</position>
<gparam>LABEL_TEXT NAND as an universal gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>102,-19</position>
<gparam>LABEL_TEXT 1.NAND AS NOT GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_TOGGLE</type>
<position>95,-24</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>102,-27.5</position>
<gparam>LABEL_TEXT 2.NAND AS AND GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>BA_NAND2</type>
<position>102,-24</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>107,-24</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>95.5,-31.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>101</ID>
<type>BA_NAND2</type>
<position>103,-32.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>95.5,-33.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>103</ID>
<type>BA_NAND2</type>
<position>112,-32.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>117.5,-32.5</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>101,-36.5</position>
<gparam>LABEL_TEXT 3.NAND AS OR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>BA_NAND2</type>
<position>97,-41.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_NAND2</type>
<position>97,-47</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>BA_NAND2</type>
<position>106,-44</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>112,-44</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>89,-41.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_TOGGLE</type>
<position>89,-47</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>141,-18.5</position>
<gparam>LABEL_TEXT 4.NAND AS NOR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>BA_NAND2</type>
<position>136,-24.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>BA_NAND2</type>
<position>136,-30</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>128,-24.5</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_TOGGLE</type>
<position>128,-30</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>118</ID>
<type>BA_NAND2</type>
<position>144,-27</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>BA_NAND2</type>
<position>152,-27</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>157,-27</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>142.5,-33.5</position>
<gparam>LABEL_TEXT 5.NAND AS XOR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>125.5,-37.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_TOGGLE</type>
<position>125,-48</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>124</ID>
<type>BA_NAND2</type>
<position>132,-42.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>BA_NAND2</type>
<position>140,-38.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>BA_NAND2</type>
<position>140,-47</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>BA_NAND2</type>
<position>149,-42.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>155,-42.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>101.5,-51.5</position>
<gparam>LABEL_TEXT 6.NAND AS XNOR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>88.5,-55.5</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>88,-66</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>133</ID>
<type>BA_NAND2</type>
<position>95,-60.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>BA_NAND2</type>
<position>103,-56.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>BA_NAND2</type>
<position>103,-65</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>BA_NAND2</type>
<position>112,-60.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>BA_NAND2</type>
<position>121,-60.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>GA_LED</type>
<position>127.5,-60.5</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>205,-9.5</position>
<gparam>LABEL_TEXT NOR as an universal gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>182,-15</position>
<gparam>LABEL_TEXT 1.NOR AS NOT GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>BE_NOR2</type>
<position>182,-21</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_TOGGLE</type>
<position>174.5,-21</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>146</ID>
<type>GA_LED</type>
<position>187.5,-21</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>226,-14</position>
<gparam>LABEL_TEXT 2.NOR AS OR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>BE_NOR2</type>
<position>211,-20.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>BE_NOR2</type>
<position>219,-20.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>225,-20.5</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>202,-19.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>202,-21.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_LABEL</type>
<position>181.5,-25.5</position>
<gparam>LABEL_TEXT 3.NOR AS AND GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>BE_NOR2</type>
<position>177,-30.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>BE_NOR2</type>
<position>177,-36.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>BE_NOR2</type>
<position>186.5,-33</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>GA_LED</type>
<position>192,-33</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_TOGGLE</type>
<position>169,-30.5</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>169,-36.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>228.5,-25</position>
<gparam>LABEL_TEXT 4.NOR AS NAND GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>BE_NOR2</type>
<position>208.5,-30.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>BE_NOR2</type>
<position>208.5,-36.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>BE_NOR2</type>
<position>218,-33</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_TOGGLE</type>
<position>200.5,-30.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>200.5,-36.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>169</ID>
<type>BE_NOR2</type>
<position>226.5,-33</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>GA_LED</type>
<position>232.5,-33</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>181.5,-41.5</position>
<gparam>LABEL_TEXT 5.NOR AS XOR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>BE_NOR2</type>
<position>171,-52</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>BE_NOR2</type>
<position>180.5,-47</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>BE_NOR2</type>
<position>180.5,-57.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>BE_NOR2</type>
<position>191,-52.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>BE_NOR2</type>
<position>202.5,-52.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>GA_LED</type>
<position>208.5,-52.5</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_TOGGLE</type>
<position>163.5,-46</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_TOGGLE</type>
<position>163.5,-58.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>228,-41.5</position>
<gparam>LABEL_TEXT 6.NOR AS XNOR GATE </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>BE_NOR2</type>
<position>220.5,-52.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>BE_NOR2</type>
<position>230,-47.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>BE_NOR2</type>
<position>230,-58</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>BE_NOR2</type>
<position>240.5,-53</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>213,-46.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>213,-59</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>192</ID>
<type>GA_LED</type>
<position>246,-53</position>
<input>
<ID>N_in0</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>298.5,-5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>272.5,-28.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>283,-28.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>315,-41.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>313.5,-52.5</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>297.5,-41</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>297.5,-47</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_AND2</type>
<position>297.5,-53.5</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_TOGGLE</type>
<position>273,-31</position>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>223</ID>
<type>AE_SMALL_INVERTER</type>
<position>276.5,-36.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_SMALL_INVERTER</type>
<position>288,-37</position>
<input>
<ID>IN_0</ID>107 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>227</ID>
<type>AE_OR2</type>
<position>308,-44</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>GA_LED</type>
<position>315,-44</position>
<input>
<ID>N_in0</ID>102 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>GA_LED</type>
<position>309,-53</position>
<input>
<ID>N_in0</ID>103 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_TOGGLE</type>
<position>283.5,-31</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_TOGGLE</type>
<position>276,-6</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_TOGGLE</type>
<position>281,-6</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>238</ID>
<type>AI_XOR2</type>
<position>295.5,-15</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>295.5,-21.5</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>GA_LED</type>
<position>302.5,-15</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>GA_LED</type>
<position>302.5,-21.5</position>
<input>
<ID>N_in0</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>276,-3</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>281,-3</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>306.5,-15</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>307,-21</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>316.5,-3.5</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>327,-3.5</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>254</ID>
<type>BA_NAND2</type>
<position>341,-14.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>BA_NAND2</type>
<position>341,-20</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>BA_NAND2</type>
<position>341,-25.5</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>BA_NAND2</type>
<position>350.5,-17</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>258</ID>
<type>BA_NAND2</type>
<position>351.5,-25.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>259</ID>
<type>GA_LED</type>
<position>356.5,-17</position>
<input>
<ID>N_in0</ID>120 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>GA_LED</type>
<position>357,-25.5</position>
<input>
<ID>N_in0</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>BA_NAND2</type>
<position>320,-9.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>BA_NAND2</type>
<position>331.5,-9.5</position>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>350.5,-7.5</position>
<gparam>LABEL_TEXT HALF ADDER WITH NAND</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>321,-31.5</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_TOGGLE</type>
<position>331.5,-31.5</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>270</ID>
<type>BE_NOR2</type>
<position>325,-37</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>BE_NOR2</type>
<position>336.5,-37</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>BE_NOR2</type>
<position>346,-43.5</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>BE_NOR2</type>
<position>346,-48.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>BE_NOR2</type>
<position>354.5,-46</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>BE_NOR2</type>
<position>363.5,-46</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>GA_LED</type>
<position>353,-54.5</position>
<input>
<ID>N_in0</ID>145 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>GA_LED</type>
<position>370,-46</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>AA_LABEL</type>
<position>357,-37</position>
<gparam>LABEL_TEXT HALF ADDER WITH NOR</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>AA_LABEL</type>
<position>405,-6.5</position>
<gparam>LABEL_TEXT HALF SUBTRACTER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>AA_AND2</type>
<position>394,-16.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AA_AND2</type>
<position>394,-22.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_TOGGLE</type>
<position>369.5,-6.5</position>
<output>
<ID>OUT_0</ID>141 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_SMALL_INVERTER</type>
<position>373,-12</position>
<input>
<ID>IN_0</ID>141 </input>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_SMALL_INVERTER</type>
<position>384.5,-12.5</position>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_OR2</type>
<position>404.5,-19.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>GA_LED</type>
<position>411.5,-19.5</position>
<input>
<ID>N_in0</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>GA_LED</type>
<position>405.5,-29</position>
<input>
<ID>N_in0</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_TOGGLE</type>
<position>380,-6.5</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_LABEL</type>
<position>394.5,-33.5</position>
<gparam>LABEL_TEXT HALF SUBTRACTER WITH NAND</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>BE_NOR2</type>
<position>346,-54.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>AA_AND2</type>
<position>394.5,-29</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>AA_TOGGLE</type>
<position>376,-36.5</position>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_TOGGLE</type>
<position>386.5,-36.5</position>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>300</ID>
<type>BA_NAND2</type>
<position>400.5,-47.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>BA_NAND2</type>
<position>400.5,-53</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>BA_NAND2</type>
<position>410,-50</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>BA_NAND2</type>
<position>411,-58.5</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>GA_LED</type>
<position>416,-50</position>
<input>
<ID>N_in0</ID>152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>305</ID>
<type>GA_LED</type>
<position>416.5,-58.5</position>
<input>
<ID>N_in0</ID>153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>306</ID>
<type>BA_NAND2</type>
<position>379.5,-42.5</position>
<input>
<ID>IN_0</ID>147 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>BA_NAND2</type>
<position>391,-42.5</position>
<input>
<ID>IN_0</ID>148 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>BA_NAND2</type>
<position>401,-58.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>AA_LABEL</type>
<position>444.5,-31.5</position>
<gparam>LABEL_TEXT HALF SUBTRACTER WITH NOR</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_TOGGLE</type>
<position>423.5,-36</position>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_TOGGLE</type>
<position>434,-36</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>312</ID>
<type>BE_NOR2</type>
<position>427.5,-41.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>BE_NOR2</type>
<position>439,-41.5</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>BE_NOR2</type>
<position>448.5,-48</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>315</ID>
<type>BE_NOR2</type>
<position>448.5,-53</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>BE_NOR2</type>
<position>457,-50.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>BE_NOR2</type>
<position>466,-50.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>GA_LED</type>
<position>455.5,-59</position>
<input>
<ID>N_in0</ID>164 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>319</ID>
<type>GA_LED</type>
<position>472.5,-50.5</position>
<input>
<ID>N_in0</ID>163 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>BE_NOR2</type>
<position>449,-59</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_TOGGLE</type>
<position>424.5,-7</position>
<output>
<ID>OUT_0</ID>165 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>322</ID>
<type>AA_TOGGLE</type>
<position>429.5,-7</position>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>323</ID>
<type>AI_XOR2</type>
<position>444,-16</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>GA_LED</type>
<position>451,-16</position>
<input>
<ID>N_in0</ID>168 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>GA_LED</type>
<position>451,-22.5</position>
<input>
<ID>N_in0</ID>169 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>443.5,-22.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>AE_SMALL_INVERTER</type>
<position>427,-11.5</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_LABEL</type>
<position>502,-5.5</position>
<gparam>LABEL_TEXT FULL ADDER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>AA_TOGGLE</type>
<position>476.5,-9.5</position>
<output>
<ID>OUT_0</ID>171 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>333</ID>
<type>AA_TOGGLE</type>
<position>481.5,-9.5</position>
<output>
<ID>OUT_0</ID>172 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_TOGGLE</type>
<position>486,-9.5</position>
<output>
<ID>OUT_0</ID>173 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_AND2</type>
<position>496.5,-20.5</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_AND2</type>
<position>496.5,-25.5</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_AND2</type>
<position>496.5,-30.5</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AI_XOR3</type>
<position>496.5,-15</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<input>
<ID>IN_2</ID>173 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>343</ID>
<type>AE_OR3</type>
<position>506,-25.5</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>175 </input>
<input>
<ID>IN_2</ID>176 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>344</ID>
<type>GA_LED</type>
<position>505.5,-15</position>
<input>
<ID>N_in0</ID>178 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>345</ID>
<type>GA_LED</type>
<position>514,-25.5</position>
<input>
<ID>N_in0</ID>177 </input>
<input>
<ID>N_in1</ID>177 </input>
<input>
<ID>N_in3</ID>177 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>AA_LABEL</type>
<position>476.5,-6.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>347</ID>
<type>AA_LABEL</type>
<position>481.5,-6.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>AA_LABEL</type>
<position>486,-6.5</position>
<gparam>LABEL_TEXT Cin</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>349</ID>
<type>AA_TOGGLE</type>
<position>477.5,-37</position>
<output>
<ID>OUT_0</ID>179 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_TOGGLE</type>
<position>485.5,-37</position>
<output>
<ID>OUT_0</ID>180 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_TOGGLE</type>
<position>493,-37</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>352</ID>
<type>BA_NAND2</type>
<position>481,-42</position>
<input>
<ID>IN_0</ID>179 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>BA_NAND2</type>
<position>489,-42</position>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>BA_NAND2</type>
<position>497,-42</position>
<input>
<ID>IN_0</ID>181 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>BA_NAND4</type>
<position>523,-60.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<input>
<ID>IN_2</ID>196 </input>
<input>
<ID>IN_3</ID>197 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>365</ID>
<type>BA_NAND4</type>
<position>524.5,-83.5</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>199 </input>
<input>
<ID>IN_2</ID>200 </input>
<input>
<ID>IN_3</ID>201 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>375</ID>
<type>BA_NAND3</type>
<position>506.5,-48.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>205 </input>
<input>
<ID>IN_2</ID>181 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>376</ID>
<type>BA_NAND3</type>
<position>506.5,-55</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>206 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>377</ID>
<type>BA_NAND3</type>
<position>506.5,-61.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>205 </input>
<input>
<ID>IN_2</ID>206 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>378</ID>
<type>BA_NAND3</type>
<position>506.5,-68.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>181 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>379</ID>
<type>BA_NAND3</type>
<position>506.5,-75</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>181 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>380</ID>
<type>BA_NAND3</type>
<position>506.5,-82.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>205 </input>
<input>
<ID>IN_2</ID>181 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>381</ID>
<type>BA_NAND3</type>
<position>506.5,-89.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>206 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>382</ID>
<type>BA_NAND3</type>
<position>506.5,-96.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>180 </input>
<input>
<ID>IN_2</ID>181 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>388</ID>
<type>GA_LED</type>
<position>530,-60.5</position>
<input>
<ID>N_in0</ID>202 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-57.5,514,-48.5</points>
<intersection>-57.5 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-57.5,520,-57.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509.5,-48.5,514,-48.5</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-18,29,-18</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509.5,-59.5,520,-59.5</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>509.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>509.5,-59.5,509.5,-55</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>-59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-20,29,-20</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509.5,-61.5,520,-61.5</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<connection>
<GID>364</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-19,37,-19</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-68.5,514,-63.5</points>
<intersection>-68.5 2</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-63.5,520,-63.5</points>
<connection>
<GID>364</GID>
<name>IN_3</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509.5,-68.5,514,-68.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-30,29.5,-30</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-80.5,514,-75</points>
<intersection>-80.5 1</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-80.5,521.5,-80.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509.5,-75,514,-75</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-32,29.5,-32</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509.5,-82.5,521.5,-82.5</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<connection>
<GID>365</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-31,37.5,-31</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509.5,-84.5,521.5,-84.5</points>
<connection>
<GID>365</GID>
<name>IN_2</name></connection>
<intersection>509.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>509.5,-89.5,509.5,-84.5</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>-84.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-39,30,-39</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>514,-96.5,514,-86.5</points>
<intersection>-96.5 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>514,-86.5,521.5,-86.5</points>
<connection>
<GID>365</GID>
<name>IN_3</name></connection>
<intersection>514 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>509.5,-96.5,514,-96.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>514 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-41,30,-41</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>526,-60.5,529,-60.5</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<connection>
<GID>388</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-40,38,-40</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<connection>
<GID>39</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527.5,-83.5,529.5,-83.5</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<connection>
<GID>390</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-48.5,30.5,-48.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>481,-73,481,-45</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<intersection>-73 5</intersection>
<intersection>-53 3</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481,-46.5,503.5,-46.5</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>481 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>481,-53,503.5,-53</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>481 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>481,-73,503.5,-73</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>481 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-50.5,30.5,-50.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>489,-82.5,489,-45</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>-82.5 5</intersection>
<intersection>-61.5 3</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>489,-48.5,503.5,-48.5</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>489 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>489,-61.5,503.5,-61.5</points>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>489 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>489,-82.5,503.5,-82.5</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>489 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-49.5,38.5,-49.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<connection>
<GID>51</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>497,-91.5,497,-45</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>-91.5 5</intersection>
<intersection>-63.5 3</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>497,-57,503.5,-57</points>
<connection>
<GID>376</GID>
<name>IN_2</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>497,-63.5,503.5,-63.5</points>
<connection>
<GID>377</GID>
<name>IN_2</name></connection>
<intersection>497 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>497,-91.5,503.5,-91.5</points>
<connection>
<GID>381</GID>
<name>IN_2</name></connection>
<intersection>497 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-18.5,58.5,-18.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-18.5,66,-18.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-27.5,62.5,-27.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-29.5,62.5,-29.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68.5,-28.5,69.5,-28.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<connection>
<GID>68</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-37,63.5,-37</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-39,63.5,-39</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-38,70.5,-38</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>79</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-25,98,-23</points>
<intersection>-25 3</intersection>
<intersection>-24 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-23,99,-23</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-24,98,-24</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>98,-25,99,-25</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>105,-24,106,-24</points>
<connection>
<GID>94</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,-31.5,100,-31.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,-33.5,100,-33.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-33.5,108,-31.5</points>
<intersection>-33.5 3</intersection>
<intersection>-32.5 4</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-31.5,109,-31.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>108,-33.5,109,-33.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>108 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106,-32.5,108,-32.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>108 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115,-32.5,116.5,-32.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>104</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-42.5,93,-40.5</points>
<intersection>-42.5 3</intersection>
<intersection>-41.5 4</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-40.5,94,-40.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>93,-42.5,94,-42.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>91,-41.5,93,-41.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-48,93,-46</points>
<intersection>-48 3</intersection>
<intersection>-47 4</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-46,94,-46</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>93,-48,94,-48</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>91,-47,93,-47</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-44,111,-44</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>109</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-43,101.5,-41.5</points>
<intersection>-43 1</intersection>
<intersection>-41.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-43,103,-43</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-41.5,101.5,-41.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-47,101.5,-45</points>
<intersection>-47 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-45,103,-45</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100,-47,101.5,-47</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-25.5,132,-23.5</points>
<intersection>-25.5 3</intersection>
<intersection>-24.5 4</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-23.5,133,-23.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,-25.5,133,-25.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-24.5,132,-24.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,-31,132,-29</points>
<intersection>-31 3</intersection>
<intersection>-30 4</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-29,133,-29</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,-31,133,-31</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>130,-30,132,-30</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-26,140,-24.5</points>
<intersection>-26 1</intersection>
<intersection>-24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,-26,141,-26</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-24.5,140,-24.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-30,140,-28</points>
<intersection>-30 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,-28,141,-28</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-30,140,-30</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-28,148,-26</points>
<intersection>-28 3</intersection>
<intersection>-27 4</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-26,149,-26</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148,-28,149,-28</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>147,-27,148,-27</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>155,-27,156,-27</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<connection>
<GID>120</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152,-42.5,154,-42.5</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,-37.5,137,-37.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>129 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>129,-41.5,129,-37.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127,-48,137,-48</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>129 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>129,-48,129,-43.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-46,136,-39.5</points>
<intersection>-46 3</intersection>
<intersection>-42.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-39.5,137,-39.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135,-42.5,136,-42.5</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136,-46,137,-46</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-41.5,144.5,-38.5</points>
<intersection>-41.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-41.5,146,-41.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-38.5,144.5,-38.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-47,144.5,-43.5</points>
<intersection>-47 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-43.5,146,-43.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-47,144.5,-47</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-55.5,100,-55.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>92 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>92,-59.5,92,-55.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-55.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-66,100,-66</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>92 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>92,-66,92,-61.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-64,99,-57.5</points>
<intersection>-64 3</intersection>
<intersection>-60.5 2</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-57.5,100,-57.5</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>98,-60.5,99,-60.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99,-64,100,-64</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-59.5,107.5,-56.5</points>
<intersection>-59.5 1</intersection>
<intersection>-56.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-59.5,109,-59.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,-56.5,107.5,-56.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107.5,-65,107.5,-61.5</points>
<intersection>-65 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-61.5,109,-61.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>107.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>106,-65,107.5,-65</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>107.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-61.5,117,-59.5</points>
<intersection>-61.5 3</intersection>
<intersection>-60.5 4</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-59.5,118,-59.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>117,-61.5,118,-61.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>115,-60.5,117,-60.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-60.5,126.5,-60.5</points>
<connection>
<GID>138</GID>
<name>N_in0</name></connection>
<connection>
<GID>137</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177.5,-22,177.5,-20</points>
<intersection>-22 3</intersection>
<intersection>-21 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177.5,-20,179,-20</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>177.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176.5,-21,177.5,-21</points>
<connection>
<GID>144</GID>
<name>OUT_0</name></connection>
<intersection>177.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>177.5,-22,179,-22</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>185,-21,186.5,-21</points>
<connection>
<GID>146</GID>
<name>N_in0</name></connection>
<connection>
<GID>142</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>216,-21.5,216,-19.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-20.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>214,-20.5,216,-20.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>216 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-19.5,208,-19.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>204,-21.5,208,-21.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-20.5,224,-20.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<connection>
<GID>151</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-31.5,173,-29.5</points>
<intersection>-31.5 3</intersection>
<intersection>-30.5 4</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,-29.5,174,-29.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>173,-31.5,174,-31.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>171,-30.5,173,-30.5</points>
<connection>
<GID>160</GID>
<name>OUT_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-37.5,173,-35.5</points>
<intersection>-37.5 3</intersection>
<intersection>-36.5 4</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>173,-35.5,174,-35.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>173,-37.5,174,-37.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>171,-36.5,173,-36.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>189.5,-33,191,-33</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<connection>
<GID>159</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-32,181.5,-30.5</points>
<intersection>-32 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-32,183.5,-32</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180,-30.5,181.5,-30.5</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-36.5,181.5,-34</points>
<intersection>-36.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-34,183.5,-34</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>181.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180,-36.5,181.5,-36.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>181.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-31.5,204.5,-29.5</points>
<intersection>-31.5 3</intersection>
<intersection>-30.5 4</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-29.5,205.5,-29.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>204.5,-31.5,205.5,-31.5</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>202.5,-30.5,204.5,-30.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204.5,-37.5,204.5,-35.5</points>
<intersection>-37.5 3</intersection>
<intersection>-36.5 4</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>204.5,-35.5,205.5,-35.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>204.5,-37.5,205.5,-37.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>204.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>202.5,-36.5,204.5,-36.5</points>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-32,213,-30.5</points>
<intersection>-32 1</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-32,215,-32</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>211.5,-30.5,213,-30.5</points>
<connection>
<GID>163</GID>
<name>OUT</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-36.5,213,-34</points>
<intersection>-36.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>213,-34,215,-34</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>211.5,-36.5,213,-36.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>213 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>222.5,-34,222.5,-32</points>
<intersection>-34 3</intersection>
<intersection>-33 4</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>222.5,-32,223.5,-32</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>222.5,-34,223.5,-34</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>222.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>221,-33,222.5,-33</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>222.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>229.5,-33,231.5,-33</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>170</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-53.5,198,-51.5</points>
<intersection>-53.5 3</intersection>
<intersection>-52.5 4</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-51.5,199.5,-51.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>198,-53.5,199.5,-53.5</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>194,-52.5,198,-52.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205.5,-52.5,207.5,-52.5</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<connection>
<GID>177</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165.5,-46,177.5,-46</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>168 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>168,-51,168,-46</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-46 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>165.5,-58.5,177.5,-58.5</points>
<connection>
<GID>181</GID>
<name>OUT_0</name></connection>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>168 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>168,-58.5,168,-53</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>-58.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-56.5,175.5,-48</points>
<intersection>-56.5 1</intersection>
<intersection>-52 2</intersection>
<intersection>-48 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-56.5,177.5,-56.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>174,-52,175.5,-52</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>175.5,-48,177.5,-48</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-51.5,185.5,-47</points>
<intersection>-51.5 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,-51.5,188,-51.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-47,185.5,-47</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185.5,-57.5,185.5,-53.5</points>
<intersection>-57.5 2</intersection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185.5,-53.5,188,-53.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>185.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-57.5,185.5,-57.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>185.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-46.5,227,-46.5</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>217.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>217.5,-51.5,217.5,-46.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-59,227,-59</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>217.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>217.5,-59,217.5,-53.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>-59 1</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>225,-57,225,-48.5</points>
<intersection>-57 1</intersection>
<intersection>-52.5 2</intersection>
<intersection>-48.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>225,-57,227,-57</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>223.5,-52.5,225,-52.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>225 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>225,-48.5,227,-48.5</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>225 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-52,235,-47.5</points>
<intersection>-52 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-52,237.5,-52</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233,-47.5,235,-47.5</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-58,235,-54</points>
<intersection>-58 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>235,-54,237.5,-54</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>233,-58,235,-58</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>243.5,-53,245,-53</points>
<connection>
<GID>192</GID>
<name>N_in0</name></connection>
<connection>
<GID>188</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-43,302.5,-41</points>
<intersection>-43 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-43,305,-43</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-41,302.5,-41</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>302.5,-47,302.5,-45</points>
<intersection>-47 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>302.5,-45,305,-45</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>302.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-47,302.5,-47</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>302.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>311,-44,314,-44</points>
<connection>
<GID>229</GID>
<name>N_in0</name></connection>
<connection>
<GID>227</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>304,-53.5,304,-53</points>
<intersection>-53.5 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>304,-53,308,-53</points>
<connection>
<GID>231</GID>
<name>N_in0</name></connection>
<intersection>304 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>300.5,-53.5,304,-53.5</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<intersection>304 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-52.5,273,-33</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 3</intersection>
<intersection>-40 1</intersection>
<intersection>-34.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>273,-40,294.5,-40</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>273,-52.5,294.5,-52.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>273,-34.5,276.5,-34.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>288,-42,288,-39</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>288,-42,294.5,-42</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>288 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276.5,-46,276.5,-38.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276.5,-46,294.5,-46</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>276.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>283.5,-54.5,283.5,-33</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-54.5 3</intersection>
<intersection>-48 1</intersection>
<intersection>-35 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>283.5,-48,294.5,-48</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>283.5,-54.5,294.5,-54.5</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>283.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>283.5,-35,288,-35</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>283.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-20.5,276,-8</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 8</intersection>
<intersection>-14 9</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>276,-20.5,292.5,-20.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>276,-14,292.5,-14</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-22.5,281,-8</points>
<connection>
<GID>236</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 3</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,-16,292.5,-16</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>281,-22.5,292.5,-22.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>281 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,-21.5,301.5,-21.5</points>
<connection>
<GID>242</GID>
<name>N_in0</name></connection>
<connection>
<GID>240</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>298.5,-15,301.5,-15</points>
<connection>
<GID>241</GID>
<name>N_in0</name></connection>
<connection>
<GID>238</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>316.5,-24.5,316.5,-5.5</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 9</intersection>
<intersection>-19 7</intersection>
<intersection>-6.5 10</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>316.5,-19,338,-19</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>316.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>316.5,-24.5,338,-24.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>316.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>316.5,-6.5,321,-6.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>316.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>327,-26.5,327,-5.5</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-26.5 9</intersection>
<intersection>-15.5 7</intersection>
<intersection>-6.5 10</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>327,-15.5,338,-15.5</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>327 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>327,-26.5,338,-26.5</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<intersection>327 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>327,-6.5,332.5,-6.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>327 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345.5,-16,345.5,-14.5</points>
<intersection>-16 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345.5,-16,347.5,-16</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>345.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>344,-14.5,345.5,-14.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<intersection>345.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>345.5,-20,345.5,-18</points>
<intersection>-20 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>345.5,-18,347.5,-18</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>345.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>344,-20,345.5,-20</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>345.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>346,-26.5,346,-24.5</points>
<intersection>-26.5 4</intersection>
<intersection>-25.5 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>346,-24.5,348.5,-24.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>346 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>344,-25.5,346,-25.5</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>346 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>346,-26.5,348.5,-26.5</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>346 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>353.5,-17,355.5,-17</points>
<connection>
<GID>259</GID>
<name>N_in0</name></connection>
<connection>
<GID>257</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>354.5,-25.5,356,-25.5</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<connection>
<GID>260</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,-21,331.5,-12.5</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>331.5,-21,338,-21</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>331.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320,-13.5,320,-12.5</points>
<connection>
<GID>262</GID>
<name>OUT</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320,-13.5,338,-13.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>320 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>321,-42.5,321,-33.5</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 8</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>321,-34,326,-34</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>321 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>321,-42.5,343,-42.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>321 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>331.5,-49.5,331.5,-33.5</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 5</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>331.5,-34,337.5,-34</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>331.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>331.5,-49.5,343,-49.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>331.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>336.5,-55.5,336.5,-40</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<intersection>-55.5 3</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>336.5,-44.5,343,-44.5</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>336.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>336.5,-55.5,343,-55.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>336.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>325,-53.5,325,-40</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>-53.5 3</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>325,-47.5,343,-47.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>325 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>325,-53.5,343,-53.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>325 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-45,350,-43.5</points>
<intersection>-45 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-45,351.5,-45</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-43.5,350,-43.5</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>350,-48.5,350,-47</points>
<intersection>-48.5 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>350,-47,351.5,-47</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>350 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>349,-48.5,350,-48.5</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>350 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>359,-47,359,-45</points>
<intersection>-47 3</intersection>
<intersection>-46 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>359,-45,360.5,-45</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>357.5,-46,359,-46</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>359 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>359,-47,360.5,-47</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>359 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>366.5,-46,369,-46</points>
<connection>
<GID>282</GID>
<name>N_in0</name></connection>
<connection>
<GID>279</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,-18.5,399,-16.5</points>
<intersection>-18.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>399,-18.5,401.5,-18.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>399 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>397,-16.5,399,-16.5</points>
<connection>
<GID>285</GID>
<name>OUT</name></connection>
<intersection>399 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>399,-22.5,399,-20.5</points>
<intersection>-22.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>399,-20.5,401.5,-20.5</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>399 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>397,-22.5,399,-22.5</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>399 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>407.5,-19.5,410.5,-19.5</points>
<connection>
<GID>292</GID>
<name>N_in0</name></connection>
<connection>
<GID>291</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>369.5,-15.5,369.5,-8.5</points>
<connection>
<GID>288</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 1</intersection>
<intersection>-10 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>369.5,-15.5,391,-15.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>369.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>369.5,-10,373,-10</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>369.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>384.5,-17.5,384.5,-14.5</points>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>384.5,-17.5,391,-17.5</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>384.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>373,-28,373,-14</points>
<connection>
<GID>289</GID>
<name>OUT_0</name></connection>
<intersection>-28 3</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>373,-21.5,391,-21.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>373 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>373,-28,391.5,-28</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>373 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>380,-30,380,-8.5</points>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection>
<intersection>-30 7</intersection>
<intersection>-23.5 1</intersection>
<intersection>-10.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>380,-23.5,391,-23.5</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>380,-10.5,384.5,-10.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>380 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>380,-30,391.5,-30</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>380 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>349,-54.5,352,-54.5</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<connection>
<GID>281</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>397.5,-29,404.5,-29</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<connection>
<GID>293</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>376,-52,376,-38.5</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>-52 7</intersection>
<intersection>-39.5 10</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>376,-52,397.5,-52</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>376 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>376,-39.5,380.5,-39.5</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>376 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>386.5,-59.5,386.5,-38.5</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>-59.5 13</intersection>
<intersection>-48.5 7</intersection>
<intersection>-39.5 10</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>386.5,-48.5,397.5,-48.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>386.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>386.5,-39.5,392,-39.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>386.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>386.5,-59.5,398,-59.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>386.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405,-49,405,-47.5</points>
<intersection>-49 1</intersection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>405,-49,407,-49</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>405 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403.5,-47.5,405,-47.5</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>405 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405,-53,405,-51</points>
<intersection>-53 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>405,-51,407,-51</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>405 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>403.5,-53,405,-53</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>405 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>405.5,-59.5,405.5,-57.5</points>
<intersection>-59.5 4</intersection>
<intersection>-58.5 5</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>405.5,-57.5,408,-57.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>405.5,-59.5,408,-59.5</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>405.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>404,-58.5,405.5,-58.5</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>413,-50,415,-50</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<connection>
<GID>304</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>414,-58.5,415.5,-58.5</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<connection>
<GID>305</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>391,-54,391,-45.5</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>391,-54,397.5,-54</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>391 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>379.5,-57.5,379.5,-45.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>-57.5 3</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>379.5,-46.5,397.5,-46.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>379.5,-57.5,398,-57.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>379.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>423.5,-47,423.5,-38</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<intersection>-47 8</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>423.5,-38.5,428.5,-38.5</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>423.5,-47,445.5,-47</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>423.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434,-60,434,-38</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<intersection>-60 8</intersection>
<intersection>-54 5</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434,-38.5,440,-38.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>434,-54,445.5,-54</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>434,-60,446,-60</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>434 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>439,-49,439,-44.5</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>439,-49,445.5,-49</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>439 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427.5,-58,427.5,-44.5</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<intersection>-58 3</intersection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427.5,-52,445.5,-52</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>427.5,-58,446,-58</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>427.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,-49.5,452.5,-48</points>
<intersection>-49.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,-49.5,454,-49.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451.5,-48,452.5,-48</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>452.5,-53,452.5,-51.5</points>
<intersection>-53 2</intersection>
<intersection>-51.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>452.5,-51.5,454,-51.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>451.5,-53,452.5,-53</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<intersection>452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>461.5,-51.5,461.5,-49.5</points>
<intersection>-51.5 3</intersection>
<intersection>-50.5 2</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>461.5,-49.5,463,-49.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>460,-50.5,461.5,-50.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>461.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>461.5,-51.5,463,-51.5</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>461.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>469,-50.5,471.5,-50.5</points>
<connection>
<GID>319</GID>
<name>N_in0</name></connection>
<connection>
<GID>317</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>452,-59,454.5,-59</points>
<connection>
<GID>318</GID>
<name>N_in0</name></connection>
<connection>
<GID>320</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>424.5,-15,424.5,-9</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>-15 9</intersection>
<intersection>-9.5 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>424.5,-15,441,-15</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>424.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>424.5,-9.5,427,-9.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>424.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>429.5,-23.5,429.5,-9</points>
<connection>
<GID>322</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 5</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>429.5,-17,441,-17</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>429.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>429.5,-23.5,440.5,-23.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>429.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>447,-16,450,-16</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<connection>
<GID>325</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>446.5,-22.5,450,-22.5</points>
<connection>
<GID>326</GID>
<name>N_in0</name></connection>
<connection>
<GID>327</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>427,-21.5,427,-13.5</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>427,-21.5,440.5,-21.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>427 0</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>476.5,-29.5,476.5,-11.5</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>-29.5 5</intersection>
<intersection>-19.5 3</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>476.5,-13,493.5,-13</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>476.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>476.5,-19.5,493.5,-19.5</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>476.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>476.5,-29.5,493.5,-29.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>476.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>481.5,-24.5,481.5,-11.5</points>
<connection>
<GID>333</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 5</intersection>
<intersection>-21.5 3</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>481.5,-15,493.5,-15</points>
<connection>
<GID>341</GID>
<name>IN_1</name></connection>
<intersection>481.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>481.5,-21.5,493.5,-21.5</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>481.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>481.5,-24.5,493.5,-24.5</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>481.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>486,-31.5,486,-11.5</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 5</intersection>
<intersection>-26.5 3</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>486,-17,493.5,-17</points>
<connection>
<GID>341</GID>
<name>IN_2</name></connection>
<intersection>486 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>486,-26.5,493.5,-26.5</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>486 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>486,-31.5,493.5,-31.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>486 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,-23.5,501,-20.5</points>
<intersection>-23.5 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>501,-23.5,503,-23.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>501 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>499.5,-20.5,501,-20.5</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>499.5,-25.5,503,-25.5</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<connection>
<GID>343</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>501,-30.5,501,-27.5</points>
<intersection>-30.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>499.5,-30.5,501,-30.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>501 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>501,-27.5,503,-27.5</points>
<connection>
<GID>343</GID>
<name>IN_2</name></connection>
<intersection>501 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>509,-25.5,515,-25.5</points>
<connection>
<GID>345</GID>
<name>N_in0</name></connection>
<connection>
<GID>345</GID>
<name>N_in1</name></connection>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<intersection>514 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>514,-25.5,514,-24.5</points>
<connection>
<GID>345</GID>
<name>N_in3</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>499.5,-15,504.5,-15</points>
<connection>
<GID>344</GID>
<name>N_in0</name></connection>
<connection>
<GID>341</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-39,482,-39</points>
<connection>
<GID>349</GID>
<name>OUT_0</name></connection>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>477.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>477.5,-94.5,477.5,-39</points>
<intersection>-94.5 12</intersection>
<intersection>-87.5 10</intersection>
<intersection>-80.5 8</intersection>
<intersection>-66.5 6</intersection>
<intersection>-59.5 4</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>477.5,-59.5,503.5,-59.5</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>477.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>477.5,-66.5,503.5,-66.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>477.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>477.5,-80.5,503.5,-80.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>477.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>477.5,-87.5,503.5,-87.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>477.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>477.5,-94.5,503.5,-94.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>477.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>485.5,-39,490,-39</points>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>485.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>485.5,-96.5,485.5,-39</points>
<intersection>-96.5 12</intersection>
<intersection>-89.5 10</intersection>
<intersection>-75 8</intersection>
<intersection>-68.5 6</intersection>
<intersection>-55 4</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>485.5,-55,503.5,-55</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<intersection>485.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>485.5,-68.5,503.5,-68.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>485.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>485.5,-75,503.5,-75</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<intersection>485.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>485.5,-89.5,503.5,-89.5</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>485.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>485.5,-96.5,503.5,-96.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>485.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>493,-39,498,-39</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>493 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>493,-98.5,493,-39</points>
<intersection>-98.5 11</intersection>
<intersection>-84.5 9</intersection>
<intersection>-77 7</intersection>
<intersection>-70.5 5</intersection>
<intersection>-50.5 3</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>493,-50.5,503.5,-50.5</points>
<connection>
<GID>375</GID>
<name>IN_2</name></connection>
<intersection>493 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>493,-70.5,503.5,-70.5</points>
<connection>
<GID>378</GID>
<name>IN_2</name></connection>
<intersection>493 2</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>493,-77,503.5,-77</points>
<connection>
<GID>379</GID>
<name>IN_2</name></connection>
<intersection>493 2</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>493,-84.5,503.5,-84.5</points>
<connection>
<GID>380</GID>
<name>IN_2</name></connection>
<intersection>493 2</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>493,-98.5,503.5,-98.5</points>
<connection>
<GID>382</GID>
<name>IN_2</name></connection>
<intersection>493 2</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,0,122.4,-60.5</PageViewport></page 9></circuit>